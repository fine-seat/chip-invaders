module chipinvaders ();
    
endmodule